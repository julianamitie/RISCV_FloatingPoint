`timescale 1ps/1ps
// 0.02 + 0.3 = 0.32
// 0_01111101_1.00110011001100110100000
// 01111101  -2
//0.01010001111010111

/* teste do módulo fpu */
module fpu_test #(parameter N = 64) ();
    
    reg clk; 
    reg rst_n;
    reg [31:0] A; 
    reg [31:0] B; 
    reg [1:0] op;
    reg start;
    wire [31:0] R;   
    wire done;    

    /* instanciação da unit under test */
    fpu uut(
        .clk(clk),
        .rst_n(rst_n),
        .A(A),
        .B(B),
        .R(R),
        .op(op),
        .start(start),
        .done(done)
    );

    /* início do testbench */
    initial begin
        clk = 0;
        rst_n = 0;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;
        
        clk = 1;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;

                clk = 0;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B", R);
        #100;

        clk = 1;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;

                clk = 0;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B", R);
        #100;

        clk = 1;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;

                clk = 0;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B", R);
        #100;

        clk = 1;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;

                clk = 0;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B", R);
        #100;

        clk = 1;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;

                clk = 0;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B", R);
        #100;

        clk = 1;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;

                clk = 0;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B", R);
        #100;

        clk = 1;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;

        clk = 0;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B", R);
        #100;

        clk = 1;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;

        clk = 0;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B", R);
        #100;

        clk = 1;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;

        clk = 0;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B", R);
        #100;

        clk = 1;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;

        clk = 0;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B", R);
        #100;

        clk = 1;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;

        clk = 0;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B", R);
        #100;

        clk = 1;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;

        clk = 0;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B", R);
        #100;

        clk = 1;
        rst_n = 1;
        A = 32'b0_01111001_01000111101100000000000;
        //0.000001010001111011  0.02 || 121 1111001
        B = 32'b0_01111101_00110011001100110100000;
        // 0.01001100110011001101  0.3  || 125 1111101
        op = 2'b00;
        start = 1;
        $monitor("R=%B \n", R);
        #100;
    
    end
endmodule