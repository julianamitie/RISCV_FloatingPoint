module rounding(
    input [22:0] fraction, 
    input [7:0] exp, 
    output reg [22:0] fractionRounded, 
    output reg [7:0] expRounded,
);

    

endmodule