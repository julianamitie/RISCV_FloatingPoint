/* descrição */
module fpu (
    input clk, rst, // clock, reset
    input [31:0] A, B, 
    output [31:0] R, 
    input [1:0] op, // operacao
    input start, 
    output done
);


endmodule